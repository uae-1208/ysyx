`include "/home/uae/ysyx/ysyx-workbench/npc/vsrc/defines.v"

module mem(
    input  wire           valid,
    input  wire           wen_mem,
    input  wire [7:0]     wmask,
    input  wire [`RegBus] waddr,
    input  wire [`RegBus] wdata,
    input  wire [2:0]     rmask,
    input  wire [`RegBus] raddr,
    output reg  [`RegBus] rdata
);
    wire           wen;
    reg  [`RegBus] rdata_temp;
    
    assign wen = wen_mem;


    import "DPI-C" function int  pmem_read(input int raddr);
    import "DPI-C" function void pmem_write(input int waddr, input int wdata, input byte wmask);
    import "DPI-C" function void ebreak(input int station, input int inst, input byte unit);


    always @(*) begin
        if(valid == 1'b1) begin // 有读写请求时
            rdata_temp = pmem_read(raddr);
            if(wen) begin // 有写请求时
                // pmem_write(waddr, 32'hdeadbeaf, wmask);
                pmem_write(waddr, wdata, wmask);
            end
        end else begin
            rdata_temp = 0;
        end
    end


    // rdata_temp -> rdata
    always @(*) begin
        case (rmask)
            `LoadBU:  rdata = {24'd0, rdata_temp[7:0]};
            `LoadHU:  rdata = {16'd0, rdata_temp[15:0]};
            // `LoadB:   rdata = {{24{rdata_temp[7]}}, rdata_temp[7:0]};
            `LoadH:   rdata = {{16{rdata_temp[15]}}, rdata_temp[15:0]};
            `LoadW:   rdata = rdata_temp;
            default:  begin
                        rdata = 0;
                        ebreak(`ABORT, 32'hdeafbeaf, `Unit_MEM);
                      end
        endcase
    end

endmodule
